library verilog;
use verilog.vl_types.all;
entity tb_ROM2 is
    generic(
        sec             : integer := 50
    );
end tb_ROM2;
