library verilog;
use verilog.vl_types.all;
entity tb_RAM1 is
    generic(
        step            : integer := 100
    );
end tb_RAM1;
