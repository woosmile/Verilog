//��� �����
module Dot_Matrix1(clk,reset,portA,portB,row,col);

//����� �����
input clk,reset;
output reg [1:0]portA,portB;
output reg [6:0]row;
output reg [4:0]col;

//ī��Ʈ ����
reg [31:0]scan_cnt;  //��ĵ �ð� ����

//portA, portB�� ��¹��� ���۷� ����
always@(posedge clk, negedge reset) begin
	if(!reset) begin
		portA <= 0;
		portB <= 0;
	end
	else begin
		portA <= 2'b01;
		portB <= 2'b01;
	end
end

//scan_cnt ���� ȸ��(�ֱ� ���� ȸ��)
always@(posedge clk, negedge reset) begin
	if(!reset) scan_cnt <= 0;
	else begin
		if(scan_cnt >= 5399999) scan_cnt <= 0;
		else scan_cnt <= scan_cnt + 1;
	end
end

//�� �ڸ� ���� ȸ��(col)
always@(posedge clk, negedge reset) begin
	if(!reset) col <= 5'b00000;
	else begin
		if(scan_cnt >= 5399999) begin
			if(col == 5'b01111) col <= 5'b11110;
			else col <= (col << 1) | 5'b00001;
		end
		else col <= col;
	end
end

//digit ���� ���� ���
always@(col) begin
	case(col)
		5'b11110 : row = 7'b1111100;
		5'b11101 : row = 7'b0010010;
		5'b11011 : row = 7'b0010001;
		5'b10111 : row = 7'b0010010;
		5'b01111 : row = 7'b1111100;
		default : row = 7'b0000000;
	endcase
end
	
endmodule
