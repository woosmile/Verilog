library verilog;
use verilog.vl_types.all;
entity tb_FSM_Moore is
    generic(
        step            : integer := 50
    );
end tb_FSM_Moore;
