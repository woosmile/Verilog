library verilog;
use verilog.vl_types.all;
entity tb_Self_Memory is
end tb_Self_Memory;
